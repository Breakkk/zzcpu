`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:45:30 11/29/2018 
// Design Name: 
// Module Name:    RegisterHeap 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RegisterHeap(

		input CLK,
		input [3:0] rdreg1_i,//A���Ĵ�����ַ
		input [3:0] rdreg2_i,//B���Ĵ�����ַ
		
		input regwrite_i,
		input [3:0] wrreg_i,//д�Ĵ�����ַ
		input [15:0] wdata_i,        //��д������
		input [15:0] epc_i,
		output [15:0] rdata1_o,
		output [15:0] rdata2_o
		
    );
	integer i;
	reg [15:0] REG_Heaps[0:15];
	initial
	begin
		for(i=15;i>=0;i=i-1)
		begin
			REG_Heaps[i] = 16'h0000;
		end
	end
	// 4'b0000 - 4'b0111: R0 - R7;
	// 4'b1000 - 4'b1011(4'b1100): SP T IH RA(EPC)
	assign rdata1_o = REG_Heaps[rdreg1_i];
	assign rdata2_o = REG_Heaps[rdreg2_i];
	
	always@(negedge CLK) begin
		if (regwrite_i) begin
			REG_Heaps[wrreg_i] <= wdata_i;
		end
		REG_Heaps[4'b1100] <= epc_i;
	end
	
	
endmodule
